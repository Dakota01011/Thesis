`timescale 1 ns / 1 ps
//////////////////////////////////////////////////////////////////////////////////
// Company: Dakota Koelling
// Engineer: Dakota Koelling
// 
// Create Date: 09/12/2016 01:49:31 PM
// Design Name: AXIS Interface
// Module Name: KNN_accelerator_v3_0_S00_AXIS
// Project Name: KNN Hardware Accelerator
// Target Devices: Zedboard, Zybo
// Tool Versions: Vivado 2016.2
// Description: 
// 
// Dependencies: 
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
//////////////////////////////////////////////////////////////////////////////////

	module KNN_accelerator_v3_0_S00_AXIS #
	(
		// AXI4Stream sink: Data Width
		parameter integer C_S_AXIS_TDATA_WIDTH	= 32
	)
	(
		// Users to add ports here
		output fifo_wren,
		output [C_S_AXIS_TDATA_WIDTH-1:0] AXIS_data,
		// User ports ends
		// Do not modify the ports beyond this line

		// AXI4Stream sink: Clock
	(* mark_debug = "true" *)	input wire  S_AXIS_ACLK,
		// AXI4Stream sink: Reset
	(* mark_debug = "true" *)	input wire  S_AXIS_ARESETN,
		// Ready to accept data in
	(* mark_debug = "true" *)	output wire  S_AXIS_TREADY,
		// Data in
	(* mark_debug = "true" *)	input wire [C_S_AXIS_TDATA_WIDTH-1 : 0] S_AXIS_TDATA,
		// Byte qualifier
	(* mark_debug = "true" *)	input wire [(C_S_AXIS_TDATA_WIDTH/8)-1 : 0] S_AXIS_TSTRB,
		// Indicates boundary of last packet
	(* mark_debug = "true" *)	input wire  S_AXIS_TLAST,
		// Data is in valid
	(* mark_debug = "true" *)	input wire  S_AXIS_TVALID
	);

	assign AXIS_data = S_AXIS_TDATA;
	assign S_AXIS_TREADY = 1;
	assign fifo_wren = S_AXIS_TVALID;

	endmodule
